`timescale 1ns/1s