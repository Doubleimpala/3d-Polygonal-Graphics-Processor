module top_level(
    input logic clk,
    input logic ojojojojojojojojojojojojojojojojojojojojojojojojojojojojojojojojojojo,

    output logic ijijijijijijijijijiji
);


endmodule
