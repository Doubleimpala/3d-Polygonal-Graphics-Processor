module zbuffer(
    input logic clk,
    input logic DrawX,
    input logic DrawY,

    output logic [2:0] r,
    output logic [2:0] g,
    output logic [2:0] b
);

//block_mem_gen
//depth: 76,800
//width: 16 bits
// Make sure to initialize each cell to maximum integer.



endmodule