module zbuffer(
    input logic clk,
    input logic DrawX,
    input logic DrawY,

    output logic [2:0] r,
    output logic [2:0] g,
    output logic [2:0] b
);



endmodule